library verilog;
use verilog.vl_types.all;
entity D_flipflop_tb is
end D_flipflop_tb;
