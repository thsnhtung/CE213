library verilog;
use verilog.vl_types.all;
entity Decoder_tb is
end Decoder_tb;
