library verilog;
use verilog.vl_types.all;
entity Mealy_tb is
end Mealy_tb;
