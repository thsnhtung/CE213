library verilog;
use verilog.vl_types.all;
entity Traffic_light_system_tb is
end Traffic_light_system_tb;
