library verilog;
use verilog.vl_types.all;
entity LoadBlock_tb is
end LoadBlock_tb;
