library verilog;
use verilog.vl_types.all;
entity registerfile_tb is
end registerfile_tb;
