library verilog;
use verilog.vl_types.all;
entity HAS_tb is
end HAS_tb;
