library verilog;
use verilog.vl_types.all;
entity DFF_tb is
end DFF_tb;
