library verilog;
use verilog.vl_types.all;
entity Decoder_1bit_tb is
end Decoder_1bit_tb;
