library verilog;
use verilog.vl_types.all;
entity Moore_tb is
end Moore_tb;
