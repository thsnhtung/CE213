library verilog;
use verilog.vl_types.all;
entity shiftReg_tb is
end shiftReg_tb;
