library verilog;
use verilog.vl_types.all;
entity D_latch_tb is
end D_latch_tb;
