library verilog;
use verilog.vl_types.all;
entity Register_1bit_tb is
end Register_1bit_tb;
