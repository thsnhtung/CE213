library verilog;
use verilog.vl_types.all;
entity Register_3bit_tb is
end Register_3bit_tb;
