library verilog;
use verilog.vl_types.all;
entity CU_tb is
end CU_tb;
