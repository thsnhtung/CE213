library verilog;
use verilog.vl_types.all;
entity StateRegiste_tb is
end StateRegiste_tb;
