module Adder_3bit (
	input [2:0]Input1,
	output wire [2:0]Result 
);
	

	assign	Result = Input1 + 1; 

endmodule

