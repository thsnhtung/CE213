library verilog;
use verilog.vl_types.all;
entity counter_1bit_tb is
end counter_1bit_tb;
