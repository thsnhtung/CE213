library verilog;
use verilog.vl_types.all;
entity Register_3bit_sync_tb is
end Register_3bit_sync_tb;
