library verilog;
use verilog.vl_types.all;
entity mealy_tb is
end mealy_tb;
