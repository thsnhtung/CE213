library verilog;
use verilog.vl_types.all;
entity register_tb is
end register_tb;
