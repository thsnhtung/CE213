library verilog;
use verilog.vl_types.all;
entity MemCell_tb is
end MemCell_tb;
