library verilog;
use verilog.vl_types.all;
entity Comparator_1bit_tb is
end Comparator_1bit_tb;
